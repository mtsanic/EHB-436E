`timescale 1ns / 1ps
module Top_Module (input A,B, output C);
AND GATE(A,B,C);
endmodule
