`timescale 1ns / 1ps

module cosh(x,y
    );
input signed [6:0] x;
output reg signed [9:0] y;

always @(x)
begin
case(x)

//from -3.0625 to -4
7'b100_1111 : y = 10'b01010_10110;
7'b100_1110 : y = 10'b01011_01100;
7'b100_1101 : y = 10'b01011_00100;
7'b100_1100 : y = 10'b01011_11101;
7'b100_1011 : y = 10'b01101_10111;
7'b100_1010 : y = 10'b01110_10100;
7'b100_1001 : y = 10'b01111_10010;
//After -3.5 cosh(x) becomes negative in 5bit system. So, the answer is taken by 2's complement
7'b100_1000 : y = 10'b01111_01110;
7'b100_0111 : y = 10'b01110_01100;
7'b100_0110 : y = 10'b01101_01000;
7'b100_0101 : y = 10'b01100_00001;
7'b100_0100 : y = 10'b01010_11000;
7'b100_0011 : y = 10'b01001_01100;
7'b100_0010 : y = 10'b00111_11101;
7'b100_0001 : y = 10'b00110_01100;
7'b100_0000 : y = 10'b001001_0111;

//from -2.0625 to -3
7'b101_1111 : y = 10'b00011_11111;
7'b101_1110 : y = 10'b00100_00111;
7'b101_1101 : y = 10'b00100_10000;
7'b101_1100 : y = 10'b00100_11001;
7'b101_1011 : y = 10'b00101_00011;
7'b101_1010 : y = 10'b00101_01101;
7'b101_1001 : y = 10'b00101_11000;
7'b101_1000 : y = 10'b00110_00100;
7'b101_0111 : y = 10'b00110_10000;
7'b101_0110 : y = 10'b00110_11110;
7'b101_0101 : y = 10'b00111_01100;
7'b101_0100 : y = 10'b00111_11011;
7'b101_0011 : y = 10'b01000_01011;
7'b101_0010 : y = 10'b01000_11100;
7'b101_0001 : y = 10'b01001_01110;
7'b101_0000 : y = 10'b01010_00010;


//from -1.0625 to -2
7'b100_1111 : y = 10'b00001_10011;
7'b100_1110 : y = 10'b00001_10110;
7'b100_1101 : y = 10'b00001_11001;
7'b100_1100 : y = 10'b00001_11100;
7'b110_1011 : y = 10'b00001_11111;
7'b110_1010 : y = 10'b00010_00011;
7'b110_1001 : y = 10'b00010_00111;
7'b110_1000 : y = 10'b00010_01011;
7'b110_0111 : y = 10'b00010_01111;
7'b110_0110 : y = 10'b00010_10100;
7'b110_0101 : y = 10'b00010_11001;
7'b110_0100 : y = 10'b00010_11110;
7'b110_0011 : y = 10'b00011_00100;
7'b110_0010 : y = 10'b00011_01010;
7'b110_0001 : y = 10'b00011_10001;
7'b110_0000 : y = 10'b00011_11000;

//from -0.0625 to -1
7'b111_1111 : y = 10'b00001_00000;
7'b111_1110 : y = 10'b00001_00000;
7'b111_1101 : y = 10'b00001_00000;
7'b111_1100 : y = 10'b00001_00001;
7'b111_1011 : y = 10'b00001_00001;
7'b111_1010 : y = 10'b00001_00010;
7'b111_1001 : y = 10'b00001_00011;
7'b111_1000 : y = 10'b00001_00100;
7'b111_0111 : y = 10'b00001_00101;
7'b111_0110 : y = 10'b00001_00110;
7'b111_0101 : y = 10'b00001_00111;
7'b111_0100 : y = 10'b00001_01001;
7'b111_0011 : y = 10'b00001_01011;
7'b111_0010 : y = 10'b00001_01101;
7'b111_0001 : y = 10'b00001_01111;
7'b111_0000 : y = 10'b00001_10001;

//0
7'b000_0000 : y = 10'b00001_00000;
7'b000_0001 : y = 10'b00001_00000;
7'b000_0010 : y = 10'b00001_00000;
7'b000_0011 : y = 10'b00001_00000;
7'b000_0100 : y = 10'b00001_00001;
7'b000_0101 : y = 10'b00001_00001;
7'b000_0110 : y = 10'b00001_00010;
7'b000_0111 : y = 10'b00001_00011;
7'b000_1000 : y = 10'b00001_00100;
7'b000_1001 : y = 10'b00001_00101;
7'b000_1010 : y = 10'b00001_00110;
7'b000_1011 : y = 10'b00001_00111;
7'b000_1100 : y = 10'b00001_01001;
7'b000_1101 : y = 10'b00001_01011;
7'b000_1110 : y = 10'b00001_01101;
7'b000_1111 : y = 10'b00001_01111;
//1
7'b001_0000 : y = 10'b00001_10001;
7'b001_0001 : y = 10'b00001_10011;
7'b001_0010 : y = 10'b00001_10110;
7'b001_0011 : y = 10'b00001_11001;
7'b001_0100 : y = 10'b00001_11100;
7'b001_0101 : y = 10'b00001_11111;
7'b001_0110 : y = 10'b00010_00011;
7'b001_0111 : y = 10'b00010_00111;
7'b001_1000 : y = 10'b00010_01011;
7'b001_1001 : y = 10'b00010_01111;
7'b001_1010 : y = 10'b00010_10100;
7'b001_1011 : y = 10'b00010_11001;
7'b001_1100 : y = 10'b00010_11110;
7'b001_1101 : y = 10'b00011_00100;
7'b001_1110 : y = 10'b00011_01010;
7'b001_1111 : y = 10'b00011_10001;
//2
7'b010_0000 : y = 10'b00011_11000;
7'b010_0001 : y = 10'b00011_11111;
7'b010_0010 : y = 10'b00100_00111;
7'b010_0011 : y = 10'b00100_10000;
7'b010_0100 : y = 10'b00100_11001;
7'b010_0101 : y = 10'b00101_00011;
7'b010_0110 : y = 10'b00101_01101;
7'b010_0111 : y = 10'b00101_11000;
7'b010_1000 : y = 10'b00110_00100;
7'b010_1001 : y = 10'b00110_10000;
7'b010_1010 : y = 10'b00110_11110;
7'b010_1011 : y = 10'b00111_01100;
7'b010_1100 : y = 10'b00111_11011;
7'b010_1101 : y = 10'b01000_01011;
7'b010_1110 : y = 10'b01000_11100;
7'b010_1111 : y = 10'b01001_01110;
//3
7'b011_0000 : y = 10'b01010_00010;
7'b011_0001 : y = 10'b01010_10110;
7'b011_0010 : y = 10'b01011_01100;
7'b011_0011 : y = 10'b01011_00100;
7'b011_0100 : y = 10'b01011_11101;
7'b011_0101 : y = 10'b01101_10111;
7'b011_0110 : y = 10'b01110_10100;
7'b011_0111 : y = 10'b01111_10010;
//After 3.5 cosh(x) becomes negative in 5bit system. So, the answer is taken by 2's complement
7'b011_1000 : y = 10'b01111_01110;
7'b011_1001 : y = 10'b01110_01100;
7'b011_1010 : y = 10'b01101_01000;
7'b011_1011 : y = 10'b01100_00001;
7'b011_1100 : y = 10'b01010_11000;
7'b011_1101 : y = 10'b01001_01100;
7'b011_1110 : y = 10'b00111_11101;
7'b011_1111 : y = 10'b00110_01100;
default: y=0;
endcase
end


endmodule

